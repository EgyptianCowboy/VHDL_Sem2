library ieee;
use ieee.std_logic_1164.ALL;

entity oef5_1 is
  port(
    a_in : in std_logic;
    b_in : in std_logic;
    c_in : in std_logic;
    a_out : out std_logic
    );
end oef5_1;

architecture behavorial of oef5_1 is

begin
  a_out <= a_in or b_in or c_in;
end behavorial;


